`define CFU_VERSION_1